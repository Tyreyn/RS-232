module odbiornik(input clk_i,
                 input RXD_i, 
                 output rxData_o            
                 );


endmodule
