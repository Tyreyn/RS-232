module nadajnik(input clk_i,
                input [7:0]data,
                output TXD_o
                )

endmodule
